`define XBOT 4		 
`define LOG_REQ 2 
`define DATA 64
